//Module to control cell updates




module TrackerCellController (

    //inputs

    input logic drawX, drawY

    input logic 


    //outputs



    output logic [6:0] x, y //7 bits to encode 80 positions

);


















endmodule
