//module for mapping user USB keycodes to their functions



//should be able to copy this from lab 5 and mofify