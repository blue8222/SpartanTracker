//Provided HDMI_Text_controller_v1_0 for HDMI AXI4 IP 
//Fall 2024 Distribution

//Modified 3/10/24 by Zuofu
//Updated 11/18/24 by Zuofu


`timescale 1 ns / 1 ps

module hdmi_text_controller_v1_0 #
(
    // Parameters of Axi Slave Bus Interface S00_AXI
    // Modify parameters as necessary for access of full VRAM range

    parameter integer C_AXI_DATA_WIDTH	= 32,
    parameter integer C_AXI_ADDR_WIDTH	= 16 // changed to 12 from 4 
)
(
    // Users to add ports here 
    
    output logic hdmi_clk_n,
    output logic hdmi_clk_p,
    output logic [2:0] hdmi_tx_n,
    output logic [2:0] hdmi_tx_p,

    // User ports ends
    // Do not modify the ports beyond this line


    // Ports of Axi Slave Bus Interface AXI
    input logic  axi_aclk,
    input logic  axi_aresetn,
    input logic [C_AXI_ADDR_WIDTH-1 : 0] axi_awaddr,
    input logic [2 : 0] axi_awprot,
    input logic  axi_awvalid,
    output logic  axi_awready,
    input logic [C_AXI_DATA_WIDTH-1 : 0] axi_wdata,
    input logic [(C_AXI_DATA_WIDTH/8)-1 : 0] axi_wstrb,
    input logic  axi_wvalid,
    output logic  axi_wready,
    output logic [1 : 0] axi_bresp,
    output logic  axi_bvalid,
    input logic  axi_bready,
    input logic [C_AXI_ADDR_WIDTH-1 : 0] axi_araddr,
    input logic [2 : 0] axi_arprot,
    input logic  axi_arvalid,
    output logic  axi_arready,
    output logic [C_AXI_DATA_WIDTH-1 : 0] axi_rdata,
    output logic [1 : 0] axi_rresp,
    output logic  axi_rvalid,
    input logic  axi_rready
);

//additional logic variables as necessary to support VGA, and HDMI modules.
    
    logic clk_25MHz, clk_125MHz;
    logic locked;
    logic [9:0] drawX;
    logic [9:0] drawY;

    logic hsync, vsync, vde;

    logic invert;
    logic [6:0] pix_code;
    logic [3:0] fg_idx;
    logic [3:0] bg_idx;
    logic [11:0] fg;
    logic [11:0] bg;
    
    logic [3:0] red, green, blue;

    // axi - vram interface
    logic axi_vram_en;
    logic [3:0] axi_vram_we;
    logic [10:0] axi_vram_addr;
    logic [31:0] axi_vram_din;
    logic [31:0] axi_vram_dout;

    // color_mapper - vram interface
    logic [10:0] cm_vram_addr;
    logic [31:0] cm_vram_dout;

    logic [9:0] cm_col, cm_row;
    logic [12:0] cm_char_ind;
    logic cm_byte_ind;

// Instantiation of Axi Bus Interface AXI
hdmi_text_controller_v1_0_AXI # ( 
    .C_S_AXI_DATA_WIDTH(C_AXI_DATA_WIDTH),
    .C_S_AXI_ADDR_WIDTH(C_AXI_ADDR_WIDTH)
) hdmi_text_controller_v1_0_AXI_inst (
    .fg_idx(fg_idx),
    .bg_idx(bg_idx),
    .fg(fg),
    .bg(bg),

    .axi_vram_en(axi_vram_en),
    .axi_vram_we(axi_vram_we),
    .axi_vram_addr(axi_vram_addr),
    .axi_vram_din(axi_vram_din),
    .axi_vram_dout(axi_vram_dout),

    .drawX(drawX),
    .drawY(drawY),
    .S_AXI_ACLK(axi_aclk),
    .S_AXI_ARESETN(axi_aresetn),
    .S_AXI_AWADDR(axi_awaddr),
    .S_AXI_AWPROT(axi_awprot),
    .S_AXI_AWVALID(axi_awvalid),
    .S_AXI_AWREADY(axi_awready),
    .S_AXI_WDATA(axi_wdata),
    .S_AXI_WSTRB(axi_wstrb),
    .S_AXI_WVALID(axi_wvalid),
    .S_AXI_WREADY(axi_wready),
    .S_AXI_BRESP(axi_bresp),
    .S_AXI_BVALID(axi_bvalid),
    .S_AXI_BREADY(axi_bready),
    .S_AXI_ARADDR(axi_araddr),
    .S_AXI_ARPROT(axi_arprot),
    .S_AXI_ARVALID(axi_arvalid),
    .S_AXI_ARREADY(axi_arready),
    .S_AXI_RDATA(axi_rdata),
    .S_AXI_RRESP(axi_rresp),
    .S_AXI_RVALID(axi_rvalid),
    .S_AXI_RREADY(axi_rready)
);


//Instiante clocking wizard, VGA sync generator modules, and VGA-HDMI IP here. For a hint, refer to the provided
//top-level from the previous lab. You should get the IP to generate a valid HDMI signal (e.g. blue screen or gradient)
//prior to working on the text drawing.

    clk_wiz_ip clk_wiz (
        .clk_out1(clk_125MHz),
        .clk_out2(clk_25MHz),
        .reset(~axi_aresetn),
        .locked(locked),
        .clk_in1(axi_aclk)
    );
    
    //VGA Sync signal generator
    vga_controller vga (
        .pixel_clk(clk_25MHz),
        .reset(~axi_aresetn),
        .hs(hsync),
        .vs(vsync),
        .active_nblank(vde),
        .drawX(drawX),
        .drawY(drawY)
    );    

    //Real Digital VGA to HDMI converter
    hdmi_tx_ip vga_to_hdmi (
        //Clocking and Reset
        .pix_clk(clk_25MHz),
        .pix_clkx5(clk_125MHz),
        .pix_clk_locked(locked),
        .rst(~axi_aresetn),

        //Color and Sync Signals
        .red(red),
        .green(green),
        .blue(blue),
        .hsync(hsync),
        .vsync(vsync),
        .vde(vde),
        
        //Differential outputs
        .TMDS_CLK_P(hdmi_clk_p),          
        .TMDS_CLK_N(hdmi_clk_n),          
        .TMDS_DATA_P(hdmi_tx_p),         
        .TMDS_DATA_N(hdmi_tx_n)          
    );

    //Color Mapper Module   
    color_mapper color_instance(
        .drawX(drawX),
        .drawY(drawY),
        .pix_code(pix_code),
        .invert(invert),
        .fg(fg),
        .bg(bg),

        .Red(red),
        .Green(green),
        .Blue(blue)
    );
    
    VRAMBlockMemory vram (
      .clka(axi_aclk),
      .ena(1'b1),
      .wea(4'b0000),
      .addra(cm_vram_addr),
      .dina(),
      .douta(cm_vram_dout),
      .clkb(axi_aclk),
      .enb(axi_vram_en),
      .web(axi_vram_we),
      .addrb(axi_vram_addr),
      .dinb(axi_vram_din),
      .doutb(axi_vram_dout)
    );

    always_comb
    begin
        cm_col = drawX / 8;
        cm_row = drawY / 16;

        cm_char_ind = (cm_row * 80) + cm_col;
        cm_vram_addr = cm_char_ind / 2;

        cm_byte_ind = cm_char_ind % 2;
        invert = cm_vram_dout[(cm_byte_ind*16)+15];
        pix_code = cm_vram_dout[(cm_byte_ind*16)+8 +: 7];
        fg_idx = cm_vram_dout[(cm_byte_ind*16)+4 +: 4];
        bg_idx = cm_vram_dout[(cm_byte_ind*16) +: 4];
    end
    
// User logic ends

endmodule
