//Module to control tracker playback




module TrackerCellController (

    //inputs

    input logic 



    //outputs



    output logic [6:0] x, y //7 bits to encode 80 positions

);


















endmodule
